magic
tech tsmc
timestamp 1754765365
<< nwell >>
rect -24 -3 61 36
rect 104 -1 151 37
<< ntransistor >>
rect -49 -18 -41 -3
rect 76 -16 84 -2
rect 125 -28 133 -14
rect -1 -42 7 -28
rect 32 -42 40 -28
<< ptransistor >>
rect -1 5 7 15
rect 32 5 40 15
rect 125 7 133 17
<< ndiffusion >>
rect -64 -4 -49 -3
rect -64 -13 -61 -4
rect -53 -13 -49 -4
rect -64 -18 -49 -13
rect -41 -4 -30 -3
rect -41 -13 -39 -4
rect -31 -13 -30 -4
rect -41 -18 -30 -13
rect 67 -3 76 -2
rect 75 -12 76 -3
rect 67 -16 76 -12
rect 84 -3 98 -2
rect 84 -12 89 -3
rect 97 -12 98 -3
rect 84 -16 98 -12
rect 113 -15 125 -14
rect 121 -24 125 -15
rect 113 -28 125 -24
rect 133 -15 143 -14
rect 133 -24 135 -15
rect 133 -28 143 -24
rect -13 -29 -1 -28
rect -5 -38 -1 -29
rect -13 -42 -1 -38
rect 7 -29 17 -28
rect 7 -38 9 -29
rect 7 -42 17 -38
rect 22 -29 32 -28
rect 30 -38 32 -29
rect 22 -42 32 -38
rect 40 -29 53 -28
rect 40 -38 44 -29
rect 52 -38 53 -29
rect 40 -42 53 -38
<< pdiffusion >>
rect -16 7 -13 15
rect -5 7 -1 15
rect -16 5 -1 7
rect 7 7 9 15
rect 7 5 17 7
rect 30 7 32 15
rect 22 5 32 7
rect 40 7 44 15
rect 52 7 53 15
rect 40 5 53 7
rect 112 9 113 17
rect 121 9 125 17
rect 112 7 125 9
rect 133 9 135 17
rect 133 7 143 9
<< ndcontact >>
rect -61 -13 -53 -4
rect -39 -13 -31 -4
rect 67 -12 75 -3
rect 89 -12 97 -3
rect 113 -24 121 -15
rect 135 -24 143 -15
rect -13 -38 -5 -29
rect 9 -38 17 -29
rect 22 -38 30 -29
rect 44 -38 52 -29
<< pdcontact >>
rect -13 7 -5 15
rect 9 7 17 15
rect 22 7 30 15
rect 44 7 52 15
rect 113 9 121 17
rect 135 9 143 17
<< psubstratepcontact >>
rect 8 -58 16 -49
rect 23 -58 31 -49
<< nsubstratencontact >>
rect 8 24 16 32
rect 23 24 31 32
rect 134 26 142 34
<< polysilicon >>
rect -49 -3 -41 37
rect -1 15 7 19
rect 32 15 40 19
rect -1 -16 7 5
rect -49 -22 -41 -18
rect -1 -28 7 -25
rect 32 -4 40 5
rect 76 -2 84 38
rect 125 17 133 21
rect 32 -28 40 -12
rect 125 -3 133 7
rect 125 -14 133 -11
rect 76 -20 84 -16
rect 125 -32 133 -28
rect -1 -46 7 -42
rect 32 -46 40 -42
<< polycontact >>
rect -53 37 -40 49
rect 75 38 84 48
rect -1 -25 7 -16
rect 32 -12 40 -4
rect 125 -11 133 -3
<< metal1 >>
rect -40 48 85 49
rect -40 38 75 48
rect 84 38 85 48
rect -40 37 85 38
rect 130 33 134 34
rect 8 32 134 33
rect 16 25 23 32
rect 16 24 17 25
rect 8 23 17 24
rect 9 15 17 23
rect 22 24 23 25
rect 31 26 134 32
rect 142 33 143 34
rect 142 26 144 33
rect 31 25 144 26
rect 22 23 31 24
rect 22 15 30 23
rect 135 17 143 25
rect -61 -4 -54 -3
rect -73 -13 -61 -4
rect -31 -5 -23 -4
rect -13 -5 -5 7
rect 44 -3 52 7
rect 113 7 121 9
rect -31 -12 32 -5
rect 44 -12 67 -3
rect 97 -8 98 -4
rect 113 -8 117 7
rect 97 -12 117 -8
rect 133 -11 158 -7
rect -73 -62 -69 -13
rect -13 -29 -5 -12
rect 44 -16 52 -12
rect 7 -25 52 -16
rect 113 -15 117 -12
rect 44 -29 52 -25
rect 9 -47 17 -38
rect 22 -47 30 -38
rect 8 -49 30 -47
rect 16 -58 23 -49
rect 135 -53 143 -24
rect 31 -58 143 -53
rect 154 -62 158 -11
rect -73 -66 158 -62
<< labels >>
rlabel metal1 -22 -8 -22 -8 1 Q
rlabel metal1 65 29 65 29 1 vdd
rlabel metal1 49 -54 49 -54 1 Gnd
rlabel metal1 -71 -11 -71 -11 3 bit
rlabel metal1 14 43 14 43 1 word
<< end >>
